//===========================================//
//  Copyright (c) Aleksandar Kostovic 2018   //
//          Matrix MAC unit package          //
//===========================================//

package mmac_pkg; //matrix-mac-package
  
 localparam DATA_WIDTH = 16; //data width of the module
  
 localparam VAR_WIDTH = 8;  //data width of internal variables
 
 localparam M_SIZE = 4; //matrix size
  
endpackage
